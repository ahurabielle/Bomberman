module mixer(input logic        active,
             input logic  [7:0] bck_r1, bck_r2,
             input logic  [7:0] bck_g1, bck_g2,
             input logic  [7:0] bck_b1, bck_b2,
             output logic [9:0] vga_r,
             output logic [9:0] vga_g,
             output logic [9:0] vga_b);

   // Vérifie qu'on est dans la zone active, sinon, c'est noir
   always @(*)
     if(active)
       begin
	  if(bck_r2 !=0)                         // on sait alors qu'on est dans le cercle blanc, donc on affiche le background2
	    begin
               vga_r <= {bck_r2, bck_r2[0], bck_r2[0]};
               vga_g <= {bck_g2, bck_g2[0], bck_g2[0]};
               vga_b <= {bck_b2, bck_b2[0], bck_b2[0]};
	    end
	  else
	    begin
	       vga_r <= {bck_r1, bck_r1[0], bck_r1[0]};
               vga_g <= {bck_g1, bck_g1[0], bck_g1[0]};
               vga_b <= {bck_b1, bck_b1[0], bck_b1[0]};
	    end // else: !if(bck_r2 !=0)
       end
     else                                     // on affiche l'autre background (sprite 1)
       {vga_r,vga_b,vga_g} <= 0;

endmodule